module DEC5T32E(I,En,Y);
    input [4:0]I;
    input En;
    output [31:0]Y;
    reg [31:0]Y;
    not i0(I_n,I);

always @(I)
    begin
        if(En==1)
            case(I)
            5'd0: Y=32'h00000001;
            5'd1: Y=32'h00000002;
            5'd2: Y=32'h00000004;
            5'd3: Y=32'h00000008;
            5'd4: Y=32'h00000010;
            5'd5: Y=32'h00000020;
            5'd6: Y=32'h00000040;
            5'd7: Y=32'h00000080;
            5'd8: Y=32'h00000100;
            5'd9: Y=32'h00000200;
            5'd10: Y=32'h00000400;
            5'd11: Y=32'h00000800;
            5'd12: Y=32'h00001000;
            5'd13: Y=32'h00002000;
            5'd14: Y=32'h00004000;
            5'd15: Y=32'h00008000;
            5'd16: Y=32'h00010000;
            5'd17: Y=32'h00020000;
            5'd18: Y=32'h00040000;
            5'd19: Y=32'h00080000;
            5'd20: Y=32'h00100000;
            5'd21: Y=32'h00200000;
            5'd22: Y=32'h00400000;
            5'd23: Y=32'h00800000;
            5'd24: Y=32'h01000000;
            5'd25: Y=32'h02000000;
            5'd26: Y=32'h04000000;
            5'd27: Y=32'h08000000;
            5'd28: Y=32'h10000000;
            5'd29: Y=32'h20000000;
            5'd30: Y=32'h40000000;
            5'd31: Y=32'h80000000;
        endcase
    else
        Y=32'd0;
    end
endmodule