module MUX32X32(
    A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    A6,
    A7,
    A8,
    A9,
    A10,
    A11,
    A12,
    A13,
    A14,
    A15,
    A16,
    A17,
    A18,
    A19,
    A20,
    A21,
    A22,
    A23,
    A24,
    A25,
    A26,
    A27,
    A28,
    A29,
    A30,
    A31,S,Y);
input [31:0]A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    A6,
    A7,
    A8,
    A9,
    A10,
    A11,
    A12,
    A13,
    A14,
    A15,
    A16,
    A17,
    A18,
    A19,
    A20,
    A21,
    A22,
    A23,
    A24,
    A25,
    A26,
    A27,
    A28,
    A29,
    A30,
    A31;
    input[4:0]S;
    output[31:0]Y;
    function[31:0]select;
    input[31:0]A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    A6,
    A7,
    A8,
    A9,
    A10,
    A11,
    A12,
    A13,
    A14,
    A15,
    A16,
    A17,
    A18,
    A19,
    A20,
    A21,
    A22,
    A23,
    A24,
    A25,
    A26,
    A27,
    A28,
    A29,
    A30,
    A31;
    input [4:0]S;
        case(S)
            5'd0:select=A0;
            5'd1:select=A1;
            5'd2:select=A2;
            5'd3:select=A3;
            5'd4:select=A4;
            5'd5:select=A5;
            5'd6:select=A6;
            5'd7:select=A7;
            5'd8:select=A8;
            5'd9:select=A9;
            5'd10:select=A10;
            5'd11:select=A11;
            5'd12:select=A12;
            5'd13:select=A13;
            5'd14:select=A14;
            5'd15:select=A15;
            5'd16:select=A16;
            5'd17:select=A17;
            5'd18:select=A18;
            5'd19:select=A19;
            5'd20:select=A20;
            5'd21:select=A21;
            5'd22:select=A22;
            5'd23:select=A23;
            5'd24:select=A24;
            5'd25:select=A25;
            5'd26:select=A26;
            5'd27:select=A27;
            5'd28:select=A28;
            5'd29:select=A29;
            5'd30:select=A30;
            5'd31:select=A31;
        endcase
    endfunction
    assign Y=select(A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    A6,
    A7,
    A8,
    A9,
    A10,
    A11,
    A12,
    A13,
    A14,
    A15,
    A16,
    A17,
    A18,
    A19,
    A20,
    A21,
    A22,
    A23,
    A24,
    A25,
    A26,
    A27,
    A28,
    A29,
    A30,
    A31,S

    );
endmodule