module MUX32X32(
    A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    A6,
    A7,
    A8,
    A9,
    A10,
    A11,
    A12,
    A13,
    A14,
    A15,
    A16,
    A17,
    A18,
    A19,
    A20,
    A21,
    A22,
    A23,
    A24,
    A25,
    A26,
    A27,
    A28,
    A29,
    A30,
    A31,S,Y);
input [31:0]A0,
    A1,
    A2,
    A3,
    A4,
    A5,
    A6,
    A7,
    A8,
    A9,
    A10,
    A11,
    A12,
    A13,
    A14,
    A15,
    A16,
    A17,
    A18,
    A19,
    A20,
    A21,
    A22,
    A23,
    A24,
    A25,
    A26,
    A27,
    A28,
    A29,
    A30,
    A31;
    input[4:0]S;
    output[31:0]Y;
    reg [31:0]Y;
    always @(S)
        begin
        case(S)
            5'd0:Y=A0;
            5'd1:Y=A1;
            5'd2:Y=A2;
            5'd3:Y=A3;
            5'd4:Y=A4;
            5'd5:Y=A5;
            5'd6:Y=A6;
            5'd7:Y=A7;
            5'd8:Y=A8;
            5'd9:Y=A9;
            5'd10:Y=A10;
            5'd11:Y=A11;
            5'd12:Y=A12;
            5'd13:Y=A13;
            5'd14:Y=A14;
            5'd15:Y=A15;
            5'd16:Y=A16;
            5'd17:Y=A17;
            5'd18:Y=A18;
            5'd19:Y=A19;
            5'd20:Y=A20;
            5'd21:Y=A21;
            5'd22:Y=A22;
            5'd23:Y=A23;
            5'd24:Y=A24;
            5'd25:Y=A25;
            5'd26:Y=A26;
            5'd27:Y=A27;
            5'd28:Y=A28;
            5'd29:Y=A29;
            5'd30:Y=A30;
            5'd31:Y=A31;
        endcase
    end
endmodule